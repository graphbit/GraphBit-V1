-----------------------------------------------------------------------
-- Character ROM that stores all all 128 ACSII characters
-- Written by Dagna Harasim, David Soofian and Charles Finkel
-----------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
entity rom_1024_8 is
port (
Clk : in std_logic;
en : in std_logic; -- Read enable
addr : in std_logic_vector(9 downto 0);
data : out std_logic_vector(7 downto 0)
);
end rom_1024_8;
architecture imp of rom_1024_8 is
type rom_type is array (0 to 1023) of std_logic_vector(7 downto 0);
constant ROM : rom_type :=
(
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",   -- 
X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
X"00", X"00", X"00", X"18", X"18", X"00", X"00", X"00",
X"10", X"38", X"7c", X"fe", X"7c", X"38", X"10", X"00",
X"38", X"7c", X"38", X"fe", X"fe", X"d6", X"10", X"38",
X"10", X"38", X"7c", X"fe", X"fe", X"7c", X"10", X"38",
X"00", X"00", X"18", X"3c", X"3c", X"18", X"00", X"00",
X"ff", X"ff", X"e7", X"c3", X"c3", X"e7", X"ff", X"ff",
X"00", X"3c", X"66", X"42", X"42", X"66", X"3c", X"00",
X"ff", X"c3", X"99", X"bd", X"bd", X"99", X"c3", X"ff",
X"0f", X"07", X"0f", X"7d", X"cc", X"cc", X"cc", X"78",
X"3c", X"66", X"66", X"66", X"3c", X"18", X"7e", X"18",
X"3f", X"33", X"3f", X"30", X"30", X"70", X"f0", X"e0",
X"7f", X"63", X"7f", X"63", X"63", X"67", X"e6", X"c0",
X"18", X"db", X"3c", X"e7", X"e7", X"3c", X"db", X"18",
X"80", X"e0", X"f8", X"fe", X"f8", X"e0", X"80", X"00",
X"02", X"0e", X"3e", X"fe", X"3e", X"0e", X"02", X"00",
X"18", X"3c", X"7e", X"18", X"18", X"7e", X"3c", X"18",
X"66", X"66", X"66", X"66", X"66", X"00", X"66", X"00",
X"7f", X"db", X"db", X"7b", X"1b", X"1b", X"1b", X"00",
X"3e", X"61", X"3c", X"66", X"66", X"3c", X"86", X"7c",
X"00", X"00", X"00", X"00", X"7e", X"7e", X"7e", X"00",
X"18", X"3c", X"7e", X"18", X"7e", X"3c", X"18", X"ff",
X"18", X"3c", X"7e", X"18", X"18", X"18", X"18", X"00",
X"18", X"18", X"18", X"18", X"7e", X"3c", X"18", X"00",
X"00", X"18", X"0c", X"fe", X"0c", X"18", X"00", X"00",
X"00", X"30", X"60", X"fe", X"60", X"30", X"00", X"00",
X"00", X"00", X"c0", X"c0", X"c0", X"fe", X"00", X"00",
X"00", X"24", X"66", X"ff", X"66", X"24", X"00", X"00",
X"00", X"18", X"3c", X"7e", X"ff", X"ff", X"00", X"00",
X"00", X"ff", X"ff", X"7e", X"3c", X"18", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",    -- 0x20 Space
X"18", X"3c", X"3c", X"18", X"18", X"00", X"18", X"00",
X"66", X"66", X"24", X"00", X"00", X"00", X"00", X"00",
X"6c", X"6c", X"fe", X"6c", X"fe", X"6c", X"6c", X"00",
X"18", X"3e", X"60", X"3c", X"06", X"7c", X"18", X"00",
X"00", X"c6", X"cc", X"18", X"30", X"66", X"c6", X"00",
X"38", X"6c", X"38", X"76", X"dc", X"cc", X"76", X"00",
X"18", X"18", X"30", X"00", X"00", X"00", X"00", X"00",
X"0c", X"18", X"30", X"30", X"30", X"18", X"0c", X"00",
X"30", X"18", X"0c", X"0c", X"0c", X"18", X"30", X"00",
X"00", X"66", X"3c", X"ff", X"3c", X"66", X"00", X"00",
X"00", X"18", X"18", X"7e", X"18", X"18", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"18", X"18", X"30",
X"00", X"00", X"00", X"7e", X"00", X"00", X"00", X"00", 
X"00", X"00", X"00", X"00", X"00", X"18", X"18", X"00",    -- 2E
X"06", X"0c", X"18", X"30", X"60", X"c0", X"80", X"00",    -- 2F
X"38", X"6c", X"c6", X"d6", X"c6", X"6c", X"38", X"00",    -- 0x30  '0'
X"18", X"38", X"18", X"18", X"18", X"18", X"7e", X"00",  
X"7c", X"c6", X"06", X"1c", X"30", X"66", X"fe", X"00",
X"7c", X"c6", X"06", X"3c", X"06", X"c6", X"7c", X"00",
X"1c", X"3c", X"6c", X"cc", X"fe", X"0c", X"1e", X"00",
X"fe", X"c0", X"c0", X"fc", X"06", X"c6", X"7c", X"00",
X"38", X"60", X"c0", X"fc", X"c6", X"c6", X"7c", X"00",
X"fe", X"c6", X"0c", X"18", X"30", X"30", X"30", X"00",
X"7c", X"c6", X"c6", X"7c", X"c6", X"c6", X"7c", X"00",
X"7c", X"c6", X"c6", X"7e", X"06", X"0c", X"78", X"00",
X"00", X"18", X"18", X"00", X"00", X"18", X"18", X"00",
X"00", X"18", X"18", X"00", X"00", X"18", X"18", X"30",
X"06", X"0c", X"18", X"30", X"18", X"0c", X"06", X"00",    -- 3C
X"00", X"00", X"7e", X"00", X"00", X"7e", X"00", X"00",    -- 3D
X"60", X"30", X"18", X"0c", X"18", X"30", X"60", X"00",    -- 3E
X"7c", X"c6", X"0c", X"18", X"18", X"00", X"18", X"00",    -- 0x3f
X"7c", X"c6", X"de", X"de", X"de", X"c0", X"78", X"00",    -- 0x40
X"38", X"6c", X"c6", X"fe", X"c6", X"c6", X"c6", X"00",    -- 0x41 'A'
X"fc", X"66", X"66", X"7c", X"66", X"66", X"fc", X"00",
X"3c", X"66", X"c0", X"c0", X"c0", X"66", X"3c", X"00",
X"f8", X"6c", X"66", X"66", X"66", X"6c", X"f8", X"00",
X"fe", X"62", X"68", X"78", X"68", X"62", X"fe", X"00",
X"fe", X"62", X"68", X"78", X"68", X"60", X"f0", X"00",
X"3c", X"66", X"c0", X"c0", X"ce", X"66", X"3a", X"00",
X"c6", X"c6", X"c6", X"fe", X"c6", X"c6", X"c6", X"00",
X"3c", X"18", X"18", X"18", X"18", X"18", X"3c", X"00",
X"1e", X"0c", X"0c", X"0c", X"cc", X"cc", X"78", X"00",
X"e6", X"66", X"6c", X"78", X"6c", X"66", X"e6", X"00",
X"f0", X"60", X"60", X"60", X"62", X"66", X"fe", X"00",
X"c6", X"ee", X"fe", X"fe", X"d6", X"c6", X"c6", X"00",
X"c6", X"e6", X"f6", X"de", X"ce", X"c6", X"c6", X"00",
X"7c", X"c6", X"c6", X"c6", X"c6", X"c6", X"7c", X"00",
X"fc", X"66", X"66", X"7c", X"60", X"60", X"f0", X"00",
X"7c", X"c6", X"c6", X"c6", X"c6", X"ce", X"7c", X"0e",
X"fc", X"66", X"66", X"7c", X"6c", X"66", X"e6", X"00",
X"3c", X"66", X"30", X"18", X"0c", X"66", X"3c", X"00",
X"7e", X"7e", X"5a", X"18", X"18", X"18", X"3c", X"00",
X"c6", X"c6", X"c6", X"c6", X"c6", X"c6", X"7c", X"00",
X"c6", X"c6", X"c6", X"c6", X"c6", X"6c", X"38", X"00",
X"c6", X"c6", X"c6", X"d6", X"d6", X"fe", X"6c", X"00",
X"c6", X"c6", X"6c", X"38", X"6c", X"c6", X"c6", X"00",
X"66", X"66", X"66", X"3c", X"18", X"18", X"3c", X"00",
X"fe", X"c6", X"8c", X"18", X"32", X"66", X"fe", X"00",
X"3c", X"30", X"30", X"30", X"30", X"30", X"3c", X"00",
X"c0", X"60", X"30", X"18", X"0c", X"06", X"02", X"00",
X"3c", X"0c", X"0c", X"0c", X"0c", X"0c", X"3c", X"00",
X"10", X"38", X"6c", X"c6", X"00", X"00", X"00", X"00",
X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"ff",
X"30", X"18", X"0c", X"00", X"00", X"00", X"00", X"00",
X"00", X"00", X"78", X"0c", X"7c", X"cc", X"76", X"00",
X"e0", X"60", X"7c", X"66", X"66", X"66", X"dc", X"00",
X"00", X"00", X"7c", X"c6", X"c0", X"c6", X"7c", X"00",
X"1c", X"0c", X"7c", X"cc", X"cc", X"cc", X"76", X"00",
X"00", X"00", X"7c", X"c6", X"fe", X"c0", X"7c", X"00",
X"3c", X"66", X"60", X"f8", X"60", X"60", X"f0", X"00",
X"00", X"00", X"76", X"cc", X"cc", X"7c", X"0c", X"f8",
X"e0", X"60", X"6c", X"76", X"66", X"66", X"e6", X"00",
X"18", X"00", X"38", X"18", X"18", X"18", X"3c", X"00",
X"06", X"00", X"06", X"06", X"06", X"66", X"66", X"3c",
X"e0", X"60", X"66", X"6c", X"78", X"6c", X"e6", X"00",
X"38", X"18", X"18", X"18", X"18", X"18", X"3c", X"00",
X"00", X"00", X"ec", X"fe", X"d6", X"d6", X"d6", X"00",
X"00", X"00", X"dc", X"66", X"66", X"66", X"66", X"00",
X"00", X"00", X"7c", X"c6", X"c6", X"c6", X"7c", X"00",
X"00", X"00", X"dc", X"66", X"66", X"7c", X"60", X"f0",
X"00", X"00", X"76", X"cc", X"cc", X"7c", X"0c", X"1e",
X"00", X"00", X"dc", X"76", X"60", X"60", X"f0", X"00",
X"00", X"00", X"7e", X"c0", X"7c", X"06", X"fc", X"00",
X"30", X"30", X"fc", X"30", X"30", X"36", X"1c", X"00",
X"00", X"00", X"cc", X"cc", X"cc", X"cc", X"76", X"00",
X"00", X"00", X"c6", X"c6", X"c6", X"6c", X"38", X"00",
X"00", X"00", X"c6", X"d6", X"d6", X"fe", X"6c", X"00",
X"00", X"00", X"c6", X"6c", X"38", X"6c", X"c6", X"00",
X"00", X"00", X"c6", X"c6", X"c6", X"7e", X"06", X"fc",
X"00", X"00", X"7e", X"4c", X"18", X"32", X"7e", X"00",
X"0e", X"18", X"18", X"70", X"18", X"18", X"0e", X"00",
X"18", X"18", X"18", X"18", X"18", X"18", X"18", X"00",
X"70", X"18", X"18", X"0e", X"18", X"18", X"70", X"00",
X"76", X"dc", X"00", X"00", X"00", X"00", X"00", X"00",
X"00", X"10", X"38", X"6c", X"c6", X"c6", X"fe", X"00"
);


begin
 process (Clk)
  begin
   if (Clk'event and Clk = '1' ) then
     if (en = '1' ) then
       data <= ROM(conv_integer(addr));
     end if;
   end if;
 end process;
end imp;